module NOT(input X,output Y);
    assign Y = ~X;
endmodule